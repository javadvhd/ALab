module Sta (
    ports
);
    
endmodule